`include "structs.sv"

module palette (
	input [2:0] palette_index,
	output RGBcolor color
);

endmodule